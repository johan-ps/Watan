1
0 0 0 0 0 g c 0 1
0 0 0 0 0 g c
0 0 0 0 0 g c
0 0 0 0 0 g c
 1 8 3 5 1 11 0 11 0 8 3 2 5 3 3 6 2 10 4 6 2 4 4 5 1 7 1 10 0 12 2 9 2 3 0 9 4 4
5
