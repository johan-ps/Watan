0
0 0 0 0 0 g c
0 0 0 0 0 g c
0 0 0 0 0 g c
0 0 0 0 0 g c
 4 7 1 10 2 5 0 8 1 4 3 9 1 11 3 10 3 6 2 4 0 9 1 3 5 11 0 2 2 5 2 3 4 12 0 8 4 6
5
